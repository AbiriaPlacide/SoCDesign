module BaudGenerator();
	
endmodule
